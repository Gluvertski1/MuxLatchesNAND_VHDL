-- Jared Day
-- 9/25/17

-- Lab 5 pt a - 2 input multiplexer with no enable line. 

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY twoinmux IS
PORT(
		i_A		:IN std_logic_vector(5 DOWNTO 0);
		o_D		:OUT std_logic_vector(7 DOWNTO 0));
END twoinmux;

ARCHITECTURE ckt of twoinmux IS
	BEGIN
		WITH i_A SELECT
		
		o_D <=	 "01111101" WHEN "000000" | "000001" | "000010" | "000011",
					 "10100011" WHEN "000100" | "000101" | "000110" | "000111",
					 "00011101" WHEN "001010" | "001011",
					 "10010010" WHEN "001000",
					 "00110000" WHEN "001001",
					 "00011101" WHEN "001110" | "001111",
					 "00010000" WHEN "001100",
					 "00110000" WHEN "001101",
					 "01111001" WHEN "010000" | "010001" | "010010" | "010011",
					 "10101110" WHEN "010100" | "010101" | "010110" | "010111",
					 "10011101" WHEN "011010" | "011011",
					 "10010110" WHEN "011000",
					 "10110000" WHEN "011001",
					 "01110111" WHEN "011100" | "011101" | "011110" | "011111",
					 "10100010" WHEN "100000" | "100001" | "100010" | "100011",
					 "10011101" WHEN "100110" | "100111",
					 "10011001" WHEN "100100",
					 "10110000" WHEN "100101",
					 "01110110"	WHEN "101000" | "101001" | "101010" | "101011",
					 "10101110" WHEN "101100" | "101101" | "101110" | "101111",
					 "10110000" WHEN "110010" | "110011",
					 "10011100" WHEN "110000", 
					 "10010000" WHEN "110001",
					 "01110101" WHEN "110100" | "110101" | "110110" | "110111",
					 "10101110" WHEN "111000" | "111001" | "111010" | "111011",
					 "10011101" WHEN "111110" | "111111",
					 "10011111" WHEN "111100",
					 "10110000" WHEN "111101",
					 "00000000" WHEN OTHERS;
END ckt;